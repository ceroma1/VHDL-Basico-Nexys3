LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY Tes0 IS
END Tes0;
 
ARCHITECTURE behavior OF Tes0 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT SupContador
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         SalidaCuenta : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';

 	--Outputs
   signal SalidaCuenta : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: SupContador PORT MAP (
          clk => clk,
          reset => reset,
          SalidaCuenta => SalidaCuenta
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 


sg_reset: process
begin		
reset<='1';
wait for 6 ns;	
reset<='0';
wait;
end process;

END;
